*Title: Case(i)

r 0 1 20
Iin 0 1 1
c 1 0 0.01 ic=0
.tran 0.02ms 20ms
.control
run
set color0 = white
plot v(1)
.endc
.end
